--
-- VHDL Architecture HEIRV32_MC.mainFSM.controller
--
-- Created:
--          by - noah.penchere.UNKNOWN (WE2330806)
--          at - 08:51:18 26.05.2023
--
-- using Mentor Graphics HDL Designer(TM) 2019.2 (Build 5)
--
ARCHITECTURE controller OF mainFSM IS
BEGIN
END ARCHITECTURE controller;

